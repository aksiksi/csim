NOR 16 51 25
NOR 16 52 26
AND 53 54 27
OR 16 55 28
OR 16 56 29
OR 16 57 30
OR 16 58 31
NOR 59 60 32
NOR 61 62 33
NOR 63 64 34
NOR 65 66 35
INV 67 36
INV 68 37
INV 69 38
INV 70 39
NAND 1 71 48
AND 1 72 49
INV 4 43
INV 5 42
INV 6 41
INV 7 40
INV 8 47
INV 9 46
INV 10 45
INV 11 44
AND 74 75 73
OR 77 78 76
INV 76 50
OR 80 81 79
OR 83 84 82
OR 86 87 85
OR 89 90 88
NAND 2 3 91
AND 76 93 92
OR 7 79 94
NAND 3 76 53
NOR 95 96 67
NOR 97 98 68
NOR 99 100 69
NOR 101 102 70
NAND 94 104 103
NOR 106 107 105
NOR 109 110 108
NOR 112 113 111
NOR 115 116 114
NOR 118 119 117
NOR 121 122 120
NOR 124 125 123
NOR 127 128 126
NOR 129 130 58
NOR 132 133 131
NOR 135 136 134
NOR 137 138 57
NOR 139 140 55
NOR 141 142 56
AND 12 143 95
AND 13 144 97
AND 14 145 99
AND 15 146 101
NOR 8 76 106
NOR 9 76 109
NOR 10 76 112
NOR 11 76 115
AND 24 73 96
AND 23 73 98
AND 22 73 100
AND 21 73 102
NOR 6 82 118
NOR 5 85 124
NOR 4 88 132
AND 92 147 61
AND 92 148 63
AND 92 149 65
AND 20 76 107
AND 19 76 110
AND 18 76 113
AND 17 76 116
NOR 4 92 139
NOR 5 92 141
NOR 6 92 137
NOR 7 92 129
AND 150 151 121
NAND 6 82 152
AND 152 153 119
AND 92 154 59
NOR 92 105 60
NOR 92 108 62
NOR 92 111 64
NOR 92 114 66
OR 156 157 155
AND 117 155 122
AND 158 159 127
NAND 5 85 160
AND 160 161 125
OR 163 164 162
AND 123 162 128
AND 92 165 130
AND 166 167 135
NAND 4 88 168
AND 168 169 133
OR 171 172 170
AND 131 170 136
AND 92 173 138
AND 92 174 140
AND 92 175 142
NAND 7 79 104
OR 177 178 176
AND 3 76 179
OR 2 179 180
AND 2 3 71
OR 182 183 181
NAND 2 179 184
NAND 176 181 51
NAND 180 184 52
NAND 82 94 185
NOR 82 94 150
NAND 85 117 186
NOR 85 117 158
NAND 88 123 187
NOR 88 123 166
NOR 2 3 74
OR 189 190 188
INV 16 54
INV 91 72
INV 1 75
INV 1 77
BUF 188 78
BUF 11 80
INV 15 81
BUF 11 83
INV 14 84
BUF 11 86
INV 13 87
BUF 11 89
INV 12 90
INV 73 93
INV 73 143
INV 73 144
INV 73 145
INV 73 146
INV 8 147
INV 9 148
INV 10 149
INV 6 151
INV 94 153
INV 103 154
INV 6 156
BUF 185 157
INV 5 159
INV 117 161
INV 5 163
BUF 186 164
INV 120 165
INV 4 167
INV 123 169
INV 4 171
BUF 187 172
INV 126 173
INV 131 174
INV 134 175
BUF 1 177
INV 91 178
INV 1 182
BUF 91 183
BUF 2 189
INV 3 190
INPUT  1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 -1
OUTPUT  25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 -1

