INV 9 5
BUF 1 12
INV 9 13
AND 12 13 7
NOR 6 14 9
NOR 3 15 11
NAND 16 17 14	
NOR 2 10 15
INV 1 18
BUF 8 19
AND 18 19 20
OR 15 20 16
OR 4 20 17
INPUT  1 2 3 4 6 8 10 -1
OUTPUT  7 9 11 5 -1
